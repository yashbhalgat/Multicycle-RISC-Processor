module RISC15_test;
	
	
endmodule